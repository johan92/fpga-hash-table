package ht_tb;

import hash_table::*;

`include "ref_hash_table.sv"
`include "ht_driver.sv"
`include "ht_monitor.sv"
`include "ht_scoreboard.sv"
`include "ht_environment.sv"

endpackage
